module simple_vectorization(output wire [3:0] out, input wire [3:0] in);
    assign out[3] = in[3];
    assign out[2] = in[2];
    assign out[1] = in[1];
    assign out[0] = in[0];
endmodule

module reverse_endianess_vectorization(output wire [3:0] out, input wire [3:0] in);
  assign out[3] = in[0];
  assign out[2] = in[1];
  assign out[1] = in[2];
  assign out[0] = in[3];
endmodule