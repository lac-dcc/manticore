// This program was cloned from: https://github.com/NYU-MLDA/OpenABC
// License: BSD 3-Clause "New" or "Revised" License

module bsg_mesh_stitch_width_p130_x_max_p2_y_max_p1
(
  outs_i,
  ins_o,
  hor_i,
  hor_o,
  ver_i,
  ver_o
);

  input [1039:0] outs_i;
  output [1039:0] ins_o;
  input [259:0] hor_i;
  output [259:0] hor_o;
  input [519:0] ver_i;
  output [519:0] ver_o;
  wire [1039:0] ins_o;
  wire [259:0] hor_o;
  wire [519:0] ver_o;
  assign ins_o[1039] = ver_i[519];
  assign ins_o[1038] = ver_i[518];
  assign ins_o[1037] = ver_i[517];
  assign ins_o[1036] = ver_i[516];
  assign ins_o[1035] = ver_i[515];
  assign ins_o[1034] = ver_i[514];
  assign ins_o[1033] = ver_i[513];
  assign ins_o[1032] = ver_i[512];
  assign ins_o[1031] = ver_i[511];
  assign ins_o[1030] = ver_i[510];
  assign ins_o[1029] = ver_i[509];
  assign ins_o[1028] = ver_i[508];
  assign ins_o[1027] = ver_i[507];
  assign ins_o[1026] = ver_i[506];
  assign ins_o[1025] = ver_i[505];
  assign ins_o[1024] = ver_i[504];
  assign ins_o[1023] = ver_i[503];
  assign ins_o[1022] = ver_i[502];
  assign ins_o[1021] = ver_i[501];
  assign ins_o[1020] = ver_i[500];
  assign ins_o[1019] = ver_i[499];
  assign ins_o[1018] = ver_i[498];
  assign ins_o[1017] = ver_i[497];
  assign ins_o[1016] = ver_i[496];
  assign ins_o[1015] = ver_i[495];
  assign ins_o[1014] = ver_i[494];
  assign ins_o[1013] = ver_i[493];
  assign ins_o[1012] = ver_i[492];
  assign ins_o[1011] = ver_i[491];
  assign ins_o[1010] = ver_i[490];
  assign ins_o[1009] = ver_i[489];
  assign ins_o[1008] = ver_i[488];
  assign ins_o[1007] = ver_i[487];
  assign ins_o[1006] = ver_i[486];
  assign ins_o[1005] = ver_i[485];
  assign ins_o[1004] = ver_i[484];
  assign ins_o[1003] = ver_i[483];
  assign ins_o[1002] = ver_i[482];
  assign ins_o[1001] = ver_i[481];
  assign ins_o[1000] = ver_i[480];
  assign ins_o[999] = ver_i[479];
  assign ins_o[998] = ver_i[478];
  assign ins_o[997] = ver_i[477];
  assign ins_o[996] = ver_i[476];
  assign ins_o[995] = ver_i[475];
  assign ins_o[994] = ver_i[474];
  assign ins_o[993] = ver_i[473];
  assign ins_o[992] = ver_i[472];
  assign ins_o[991] = ver_i[471];
  assign ins_o[990] = ver_i[470];
  assign ins_o[989] = ver_i[469];
  assign ins_o[988] = ver_i[468];
  assign ins_o[987] = ver_i[467];
  assign ins_o[986] = ver_i[466];
  assign ins_o[985] = ver_i[465];
  assign ins_o[984] = ver_i[464];
  assign ins_o[983] = ver_i[463];
  assign ins_o[982] = ver_i[462];
  assign ins_o[981] = ver_i[461];
  assign ins_o[980] = ver_i[460];
  assign ins_o[979] = ver_i[459];
  assign ins_o[978] = ver_i[458];
  assign ins_o[977] = ver_i[457];
  assign ins_o[976] = ver_i[456];
  assign ins_o[975] = ver_i[455];
  assign ins_o[974] = ver_i[454];
  assign ins_o[973] = ver_i[453];
  assign ins_o[972] = ver_i[452];
  assign ins_o[971] = ver_i[451];
  assign ins_o[970] = ver_i[450];
  assign ins_o[969] = ver_i[449];
  assign ins_o[968] = ver_i[448];
  assign ins_o[967] = ver_i[447];
  assign ins_o[966] = ver_i[446];
  assign ins_o[965] = ver_i[445];
  assign ins_o[964] = ver_i[444];
  assign ins_o[963] = ver_i[443];
  assign ins_o[962] = ver_i[442];
  assign ins_o[961] = ver_i[441];
  assign ins_o[960] = ver_i[440];
  assign ins_o[959] = ver_i[439];
  assign ins_o[958] = ver_i[438];
  assign ins_o[957] = ver_i[437];
  assign ins_o[956] = ver_i[436];
  assign ins_o[955] = ver_i[435];
  assign ins_o[954] = ver_i[434];
  assign ins_o[953] = ver_i[433];
  assign ins_o[952] = ver_i[432];
  assign ins_o[951] = ver_i[431];
  assign ins_o[950] = ver_i[430];
  assign ins_o[949] = ver_i[429];
  assign ins_o[948] = ver_i[428];
  assign ins_o[947] = ver_i[427];
  assign ins_o[946] = ver_i[426];
  assign ins_o[945] = ver_i[425];
  assign ins_o[944] = ver_i[424];
  assign ins_o[943] = ver_i[423];
  assign ins_o[942] = ver_i[422];
  assign ins_o[941] = ver_i[421];
  assign ins_o[940] = ver_i[420];
  assign ins_o[939] = ver_i[419];
  assign ins_o[938] = ver_i[418];
  assign ins_o[937] = ver_i[417];
  assign ins_o[936] = ver_i[416];
  assign ins_o[935] = ver_i[415];
  assign ins_o[934] = ver_i[414];
  assign ins_o[933] = ver_i[413];
  assign ins_o[932] = ver_i[412];
  assign ins_o[931] = ver_i[411];
  assign ins_o[930] = ver_i[410];
  assign ins_o[929] = ver_i[409];
  assign ins_o[928] = ver_i[408];
  assign ins_o[927] = ver_i[407];
  assign ins_o[926] = ver_i[406];
  assign ins_o[925] = ver_i[405];
  assign ins_o[924] = ver_i[404];
  assign ins_o[923] = ver_i[403];
  assign ins_o[922] = ver_i[402];
  assign ins_o[921] = ver_i[401];
  assign ins_o[920] = ver_i[400];
  assign ins_o[919] = ver_i[399];
  assign ins_o[918] = ver_i[398];
  assign ins_o[917] = ver_i[397];
  assign ins_o[916] = ver_i[396];
  assign ins_o[915] = ver_i[395];
  assign ins_o[914] = ver_i[394];
  assign ins_o[913] = ver_i[393];
  assign ins_o[912] = ver_i[392];
  assign ins_o[911] = ver_i[391];
  assign ins_o[910] = ver_i[390];
  assign ins_o[909] = ver_i[259];
  assign ins_o[908] = ver_i[258];
  assign ins_o[907] = ver_i[257];
  assign ins_o[906] = ver_i[256];
  assign ins_o[905] = ver_i[255];
  assign ins_o[904] = ver_i[254];
  assign ins_o[903] = ver_i[253];
  assign ins_o[902] = ver_i[252];
  assign ins_o[901] = ver_i[251];
  assign ins_o[900] = ver_i[250];
  assign ins_o[899] = ver_i[249];
  assign ins_o[898] = ver_i[248];
  assign ins_o[897] = ver_i[247];
  assign ins_o[896] = ver_i[246];
  assign ins_o[895] = ver_i[245];
  assign ins_o[894] = ver_i[244];
  assign ins_o[893] = ver_i[243];
  assign ins_o[892] = ver_i[242];
  assign ins_o[891] = ver_i[241];
  assign ins_o[890] = ver_i[240];
  assign ins_o[889] = ver_i[239];
  assign ins_o[888] = ver_i[238];
  assign ins_o[887] = ver_i[237];
  assign ins_o[886] = ver_i[236];
  assign ins_o[885] = ver_i[235];
  assign ins_o[884] = ver_i[234];
  assign ins_o[883] = ver_i[233];
  assign ins_o[882] = ver_i[232];
  assign ins_o[881] = ver_i[231];
  assign ins_o[880] = ver_i[230];
  assign ins_o[879] = ver_i[229];
  assign ins_o[878] = ver_i[228];
  assign ins_o[877] = ver_i[227];
  assign ins_o[876] = ver_i[226];
  assign ins_o[875] = ver_i[225];
  assign ins_o[874] = ver_i[224];
  assign ins_o[873] = ver_i[223];
  assign ins_o[872] = ver_i[222];
  assign ins_o[871] = ver_i[221];
  assign ins_o[870] = ver_i[220];
  assign ins_o[869] = ver_i[219];
  assign ins_o[868] = ver_i[218];
  assign ins_o[867] = ver_i[217];
  assign ins_o[866] = ver_i[216];
  assign ins_o[865] = ver_i[215];
  assign ins_o[864] = ver_i[214];
  assign ins_o[863] = ver_i[213];
  assign ins_o[862] = ver_i[212];
  assign ins_o[861] = ver_i[211];
  assign ins_o[860] = ver_i[210];
  assign ins_o[859] = ver_i[209];
  assign ins_o[858] = ver_i[208];
  assign ins_o[857] = ver_i[207];
  assign ins_o[856] = ver_i[206];
  assign ins_o[855] = ver_i[205];
  assign ins_o[854] = ver_i[204];
  assign ins_o[853] = ver_i[203];
  assign ins_o[852] = ver_i[202];
  assign ins_o[851] = ver_i[201];
  assign ins_o[850] = ver_i[200];
  assign ins_o[849] = ver_i[199];
  assign ins_o[848] = ver_i[198];
  assign ins_o[847] = ver_i[197];
  assign ins_o[846] = ver_i[196];
  assign ins_o[845] = ver_i[195];
  assign ins_o[844] = ver_i[194];
  assign ins_o[843] = ver_i[193];
  assign ins_o[842] = ver_i[192];
  assign ins_o[841] = ver_i[191];
  assign ins_o[840] = ver_i[190];
  assign ins_o[839] = ver_i[189];
  assign ins_o[838] = ver_i[188];
  assign ins_o[837] = ver_i[187];
  assign ins_o[836] = ver_i[186];
  assign ins_o[835] = ver_i[185];
  assign ins_o[834] = ver_i[184];
  assign ins_o[833] = ver_i[183];
  assign ins_o[832] = ver_i[182];
  assign ins_o[831] = ver_i[181];
  assign ins_o[830] = ver_i[180];
  assign ins_o[829] = ver_i[179];
  assign ins_o[828] = ver_i[178];
  assign ins_o[827] = ver_i[177];
  assign ins_o[826] = ver_i[176];
  assign ins_o[825] = ver_i[175];
  assign ins_o[824] = ver_i[174];
  assign ins_o[823] = ver_i[173];
  assign ins_o[822] = ver_i[172];
  assign ins_o[821] = ver_i[171];
  assign ins_o[820] = ver_i[170];
  assign ins_o[819] = ver_i[169];
  assign ins_o[818] = ver_i[168];
  assign ins_o[817] = ver_i[167];
  assign ins_o[816] = ver_i[166];
  assign ins_o[815] = ver_i[165];
  assign ins_o[814] = ver_i[164];
  assign ins_o[813] = ver_i[163];
  assign ins_o[812] = ver_i[162];
  assign ins_o[811] = ver_i[161];
  assign ins_o[810] = ver_i[160];
  assign ins_o[809] = ver_i[159];
  assign ins_o[808] = ver_i[158];
  assign ins_o[807] = ver_i[157];
  assign ins_o[806] = ver_i[156];
  assign ins_o[805] = ver_i[155];
  assign ins_o[804] = ver_i[154];
  assign ins_o[803] = ver_i[153];
  assign ins_o[802] = ver_i[152];
  assign ins_o[801] = ver_i[151];
  assign ins_o[800] = ver_i[150];
  assign ins_o[799] = ver_i[149];
  assign ins_o[798] = ver_i[148];
  assign ins_o[797] = ver_i[147];
  assign ins_o[796] = ver_i[146];
  assign ins_o[795] = ver_i[145];
  assign ins_o[794] = ver_i[144];
  assign ins_o[793] = ver_i[143];
  assign ins_o[792] = ver_i[142];
  assign ins_o[791] = ver_i[141];
  assign ins_o[790] = ver_i[140];
  assign ins_o[789] = ver_i[139];
  assign ins_o[788] = ver_i[138];
  assign ins_o[787] = ver_i[137];
  assign ins_o[786] = ver_i[136];
  assign ins_o[785] = ver_i[135];
  assign ins_o[784] = ver_i[134];
  assign ins_o[783] = ver_i[133];
  assign ins_o[782] = ver_i[132];
  assign ins_o[781] = ver_i[131];
  assign ins_o[780] = ver_i[130];
  assign ins_o[779] = hor_i[259];
  assign ins_o[778] = hor_i[258];
  assign ins_o[777] = hor_i[257];
  assign ins_o[776] = hor_i[256];
  assign ins_o[775] = hor_i[255];
  assign ins_o[774] = hor_i[254];
  assign ins_o[773] = hor_i[253];
  assign ins_o[772] = hor_i[252];
  assign ins_o[771] = hor_i[251];
  assign ins_o[770] = hor_i[250];
  assign ins_o[769] = hor_i[249];
  assign ins_o[768] = hor_i[248];
  assign ins_o[767] = hor_i[247];
  assign ins_o[766] = hor_i[246];
  assign ins_o[765] = hor_i[245];
  assign ins_o[764] = hor_i[244];
  assign ins_o[763] = hor_i[243];
  assign ins_o[762] = hor_i[242];
  assign ins_o[761] = hor_i[241];
  assign ins_o[760] = hor_i[240];
  assign ins_o[759] = hor_i[239];
  assign ins_o[758] = hor_i[238];
  assign ins_o[757] = hor_i[237];
  assign ins_o[756] = hor_i[236];
  assign ins_o[755] = hor_i[235];
  assign ins_o[754] = hor_i[234];
  assign ins_o[753] = hor_i[233];
  assign ins_o[752] = hor_i[232];
  assign ins_o[751] = hor_i[231];
  assign ins_o[750] = hor_i[230];
  assign ins_o[749] = hor_i[229];
  assign ins_o[748] = hor_i[228];
  assign ins_o[747] = hor_i[227];
  assign ins_o[746] = hor_i[226];
  assign ins_o[745] = hor_i[225];
  assign ins_o[744] = hor_i[224];
  assign ins_o[743] = hor_i[223];
  assign ins_o[742] = hor_i[222];
  assign ins_o[741] = hor_i[221];
  assign ins_o[740] = hor_i[220];
  assign ins_o[739] = hor_i[219];
  assign ins_o[738] = hor_i[218];
  assign ins_o[737] = hor_i[217];
  assign ins_o[736] = hor_i[216];
  assign ins_o[735] = hor_i[215];
  assign ins_o[734] = hor_i[214];
  assign ins_o[733] = hor_i[213];
  assign ins_o[732] = hor_i[212];
  assign ins_o[731] = hor_i[211];
  assign ins_o[730] = hor_i[210];
  assign ins_o[729] = hor_i[209];
  assign ins_o[728] = hor_i[208];
  assign ins_o[727] = hor_i[207];
  assign ins_o[726] = hor_i[206];
  assign ins_o[725] = hor_i[205];
  assign ins_o[724] = hor_i[204];
  assign ins_o[723] = hor_i[203];
  assign ins_o[722] = hor_i[202];
  assign ins_o[721] = hor_i[201];
  assign ins_o[720] = hor_i[200];
  assign ins_o[719] = hor_i[199];
  assign ins_o[718] = hor_i[198];
  assign ins_o[717] = hor_i[197];
  assign ins_o[716] = hor_i[196];
  assign ins_o[715] = hor_i[195];
  assign ins_o[714] = hor_i[194];
  assign ins_o[713] = hor_i[193];
  assign ins_o[712] = hor_i[192];
  assign ins_o[711] = hor_i[191];
  assign ins_o[710] = hor_i[190];
  assign ins_o[709] = hor_i[189];
  assign ins_o[708] = hor_i[188];
  assign ins_o[707] = hor_i[187];
  assign ins_o[706] = hor_i[186];
  assign ins_o[705] = hor_i[185];
  assign ins_o[704] = hor_i[184];
  assign ins_o[703] = hor_i[183];
  assign ins_o[702] = hor_i[182];
  assign ins_o[701] = hor_i[181];
  assign ins_o[700] = hor_i[180];
  assign ins_o[699] = hor_i[179];
  assign ins_o[698] = hor_i[178];
  assign ins_o[697] = hor_i[177];
  assign ins_o[696] = hor_i[176];
  assign ins_o[695] = hor_i[175];
  assign ins_o[694] = hor_i[174];
  assign ins_o[693] = hor_i[173];
  assign ins_o[692] = hor_i[172];
  assign ins_o[691] = hor_i[171];
  assign ins_o[690] = hor_i[170];
  assign ins_o[689] = hor_i[169];
  assign ins_o[688] = hor_i[168];
  assign ins_o[687] = hor_i[167];
  assign ins_o[686] = hor_i[166];
  assign ins_o[685] = hor_i[165];
  assign ins_o[684] = hor_i[164];
  assign ins_o[683] = hor_i[163];
  assign ins_o[682] = hor_i[162];
  assign ins_o[681] = hor_i[161];
  assign ins_o[680] = hor_i[160];
  assign ins_o[679] = hor_i[159];
  assign ins_o[678] = hor_i[158];
  assign ins_o[677] = hor_i[157];
  assign ins_o[676] = hor_i[156];
  assign ins_o[675] = hor_i[155];
  assign ins_o[674] = hor_i[154];
  assign ins_o[673] = hor_i[153];
  assign ins_o[672] = hor_i[152];
  assign ins_o[671] = hor_i[151];
  assign ins_o[670] = hor_i[150];
  assign ins_o[669] = hor_i[149];
  assign ins_o[668] = hor_i[148];
  assign ins_o[667] = hor_i[147];
  assign ins_o[666] = hor_i[146];
  assign ins_o[665] = hor_i[145];
  assign ins_o[664] = hor_i[144];
  assign ins_o[663] = hor_i[143];
  assign ins_o[662] = hor_i[142];
  assign ins_o[661] = hor_i[141];
  assign ins_o[660] = hor_i[140];
  assign ins_o[659] = hor_i[139];
  assign ins_o[658] = hor_i[138];
  assign ins_o[657] = hor_i[137];
  assign ins_o[656] = hor_i[136];
  assign ins_o[655] = hor_i[135];
  assign ins_o[654] = hor_i[134];
  assign ins_o[653] = hor_i[133];
  assign ins_o[652] = hor_i[132];
  assign ins_o[651] = hor_i[131];
  assign ins_o[650] = hor_i[130];
  assign ins_o[649] = outs_i[259];
  assign ins_o[648] = outs_i[258];
  assign ins_o[647] = outs_i[257];
  assign ins_o[646] = outs_i[256];
  assign ins_o[645] = outs_i[255];
  assign ins_o[644] = outs_i[254];
  assign ins_o[643] = outs_i[253];
  assign ins_o[642] = outs_i[252];
  assign ins_o[641] = outs_i[251];
  assign ins_o[640] = outs_i[250];
  assign ins_o[639] = outs_i[249];
  assign ins_o[638] = outs_i[248];
  assign ins_o[637] = outs_i[247];
  assign ins_o[636] = outs_i[246];
  assign ins_o[635] = outs_i[245];
  assign ins_o[634] = outs_i[244];
  assign ins_o[633] = outs_i[243];
  assign ins_o[632] = outs_i[242];
  assign ins_o[631] = outs_i[241];
  assign ins_o[630] = outs_i[240];
  assign ins_o[629] = outs_i[239];
  assign ins_o[628] = outs_i[238];
  assign ins_o[627] = outs_i[237];
  assign ins_o[626] = outs_i[236];
  assign ins_o[625] = outs_i[235];
  assign ins_o[624] = outs_i[234];
  assign ins_o[623] = outs_i[233];
  assign ins_o[622] = outs_i[232];
  assign ins_o[621] = outs_i[231];
  assign ins_o[620] = outs_i[230];
  assign ins_o[619] = outs_i[229];
  assign ins_o[618] = outs_i[228];
  assign ins_o[617] = outs_i[227];
  assign ins_o[616] = outs_i[226];
  assign ins_o[615] = outs_i[225];
  assign ins_o[614] = outs_i[224];
  assign ins_o[613] = outs_i[223];
  assign ins_o[612] = outs_i[222];
  assign ins_o[611] = outs_i[221];
  assign ins_o[610] = outs_i[220];
  assign ins_o[609] = outs_i[219];
  assign ins_o[608] = outs_i[218];
  assign ins_o[607] = outs_i[217];
  assign ins_o[606] = outs_i[216];
  assign ins_o[605] = outs_i[215];
  assign ins_o[604] = outs_i[214];
  assign ins_o[603] = outs_i[213];
  assign ins_o[602] = outs_i[212];
  assign ins_o[601] = outs_i[211];
  assign ins_o[600] = outs_i[210];
  assign ins_o[599] = outs_i[209];
  assign ins_o[598] = outs_i[208];
  assign ins_o[597] = outs_i[207];
  assign ins_o[596] = outs_i[206];
  assign ins_o[595] = outs_i[205];
  assign ins_o[594] = outs_i[204];
  assign ins_o[593] = outs_i[203];
  assign ins_o[592] = outs_i[202];
  assign ins_o[591] = outs_i[201];
  assign ins_o[590] = outs_i[200];
  assign ins_o[589] = outs_i[199];
  assign ins_o[588] = outs_i[198];
  assign ins_o[587] = outs_i[197];
  assign ins_o[586] = outs_i[196];
  assign ins_o[585] = outs_i[195];
  assign ins_o[584] = outs_i[194];
  assign ins_o[583] = outs_i[193];
  assign ins_o[582] = outs_i[192];
  assign ins_o[581] = outs_i[191];
  assign ins_o[580] = outs_i[190];
  assign ins_o[579] = outs_i[189];
  assign ins_o[578] = outs_i[188];
  assign ins_o[577] = outs_i[187];
  assign ins_o[576] = outs_i[186];
  assign ins_o[575] = outs_i[185];
  assign ins_o[574] = outs_i[184];
  assign ins_o[573] = outs_i[183];
  assign ins_o[572] = outs_i[182];
  assign ins_o[571] = outs_i[181];
  assign ins_o[570] = outs_i[180];
  assign ins_o[569] = outs_i[179];
  assign ins_o[568] = outs_i[178];
  assign ins_o[567] = outs_i[177];
  assign ins_o[566] = outs_i[176];
  assign ins_o[565] = outs_i[175];
  assign ins_o[564] = outs_i[174];
  assign ins_o[563] = outs_i[173];
  assign ins_o[562] = outs_i[172];
  assign ins_o[561] = outs_i[171];
  assign ins_o[560] = outs_i[170];
  assign ins_o[559] = outs_i[169];
  assign ins_o[558] = outs_i[168];
  assign ins_o[557] = outs_i[167];
  assign ins_o[556] = outs_i[166];
  assign ins_o[555] = outs_i[165];
  assign ins_o[554] = outs_i[164];
  assign ins_o[553] = outs_i[163];
  assign ins_o[552] = outs_i[162];
  assign ins_o[551] = outs_i[161];
  assign ins_o[550] = outs_i[160];
  assign ins_o[549] = outs_i[159];
  assign ins_o[548] = outs_i[158];
  assign ins_o[547] = outs_i[157];
  assign ins_o[546] = outs_i[156];
  assign ins_o[545] = outs_i[155];
  assign ins_o[544] = outs_i[154];
  assign ins_o[543] = outs_i[153];
  assign ins_o[542] = outs_i[152];
  assign ins_o[541] = outs_i[151];
  assign ins_o[540] = outs_i[150];
  assign ins_o[539] = outs_i[149];
  assign ins_o[538] = outs_i[148];
  assign ins_o[537] = outs_i[147];
  assign ins_o[536] = outs_i[146];
  assign ins_o[535] = outs_i[145];
  assign ins_o[534] = outs_i[144];
  assign ins_o[533] = outs_i[143];
  assign ins_o[532] = outs_i[142];
  assign ins_o[531] = outs_i[141];
  assign ins_o[530] = outs_i[140];
  assign ins_o[529] = outs_i[139];
  assign ins_o[528] = outs_i[138];
  assign ins_o[527] = outs_i[137];
  assign ins_o[526] = outs_i[136];
  assign ins_o[525] = outs_i[135];
  assign ins_o[524] = outs_i[134];
  assign ins_o[523] = outs_i[133];
  assign ins_o[522] = outs_i[132];
  assign ins_o[521] = outs_i[131];
  assign ins_o[520] = outs_i[130];
  assign ins_o[519] = ver_i[389];
  assign ins_o[518] = ver_i[388];
  assign ins_o[517] = ver_i[387];
  assign ins_o[516] = ver_i[386];
  assign ins_o[515] = ver_i[385];
  assign ins_o[514] = ver_i[384];
  assign ins_o[513] = ver_i[383];
  assign ins_o[512] = ver_i[382];
  assign ins_o[511] = ver_i[381];
  assign ins_o[510] = ver_i[380];
  assign ins_o[509] = ver_i[379];
  assign ins_o[508] = ver_i[378];
  assign ins_o[507] = ver_i[377];
  assign ins_o[506] = ver_i[376];
  assign ins_o[505] = ver_i[375];
  assign ins_o[504] = ver_i[374];
  assign ins_o[503] = ver_i[373];
  assign ins_o[502] = ver_i[372];
  assign ins_o[501] = ver_i[371];
  assign ins_o[500] = ver_i[370];
  assign ins_o[499] = ver_i[369];
  assign ins_o[498] = ver_i[368];
  assign ins_o[497] = ver_i[367];
  assign ins_o[496] = ver_i[366];
  assign ins_o[495] = ver_i[365];
  assign ins_o[494] = ver_i[364];
  assign ins_o[493] = ver_i[363];
  assign ins_o[492] = ver_i[362];
  assign ins_o[491] = ver_i[361];
  assign ins_o[490] = ver_i[360];
  assign ins_o[489] = ver_i[359];
  assign ins_o[488] = ver_i[358];
  assign ins_o[487] = ver_i[357];
  assign ins_o[486] = ver_i[356];
  assign ins_o[485] = ver_i[355];
  assign ins_o[484] = ver_i[354];
  assign ins_o[483] = ver_i[353];
  assign ins_o[482] = ver_i[352];
  assign ins_o[481] = ver_i[351];
  assign ins_o[480] = ver_i[350];
  assign ins_o[479] = ver_i[349];
  assign ins_o[478] = ver_i[348];
  assign ins_o[477] = ver_i[347];
  assign ins_o[476] = ver_i[346];
  assign ins_o[475] = ver_i[345];
  assign ins_o[474] = ver_i[344];
  assign ins_o[473] = ver_i[343];
  assign ins_o[472] = ver_i[342];
  assign ins_o[471] = ver_i[341];
  assign ins_o[470] = ver_i[340];
  assign ins_o[469] = ver_i[339];
  assign ins_o[468] = ver_i[338];
  assign ins_o[467] = ver_i[337];
  assign ins_o[466] = ver_i[336];
  assign ins_o[465] = ver_i[335];
  assign ins_o[464] = ver_i[334];
  assign ins_o[463] = ver_i[333];
  assign ins_o[462] = ver_i[332];
  assign ins_o[461] = ver_i[331];
  assign ins_o[460] = ver_i[330];
  assign ins_o[459] = ver_i[329];
  assign ins_o[458] = ver_i[328];
  assign ins_o[457] = ver_i[327];
  assign ins_o[456] = ver_i[326];
  assign ins_o[455] = ver_i[325];
  assign ins_o[454] = ver_i[324];
  assign ins_o[453] = ver_i[323];
  assign ins_o[452] = ver_i[322];
  assign ins_o[451] = ver_i[321];
  assign ins_o[450] = ver_i[320];
  assign ins_o[449] = ver_i[319];
  assign ins_o[448] = ver_i[318];
  assign ins_o[447] = ver_i[317];
  assign ins_o[446] = ver_i[316];
  assign ins_o[445] = ver_i[315];
  assign ins_o[444] = ver_i[314];
  assign ins_o[443] = ver_i[313];
  assign ins_o[442] = ver_i[312];
  assign ins_o[441] = ver_i[311];
  assign ins_o[440] = ver_i[310];
  assign ins_o[439] = ver_i[309];
  assign ins_o[438] = ver_i[308];
  assign ins_o[437] = ver_i[307];
  assign ins_o[436] = ver_i[306];
  assign ins_o[435] = ver_i[305];
  assign ins_o[434] = ver_i[304];
  assign ins_o[433] = ver_i[303];
  assign ins_o[432] = ver_i[302];
  assign ins_o[431] = ver_i[301];
  assign ins_o[430] = ver_i[300];
  assign ins_o[429] = ver_i[299];
  assign ins_o[428] = ver_i[298];
  assign ins_o[427] = ver_i[297];
  assign ins_o[426] = ver_i[296];
  assign ins_o[425] = ver_i[295];
  assign ins_o[424] = ver_i[294];
  assign ins_o[423] = ver_i[293];
  assign ins_o[422] = ver_i[292];
  assign ins_o[421] = ver_i[291];
  assign ins_o[420] = ver_i[290];
  assign ins_o[419] = ver_i[289];
  assign ins_o[418] = ver_i[288];
  assign ins_o[417] = ver_i[287];
  assign ins_o[416] = ver_i[286];
  assign ins_o[415] = ver_i[285];
  assign ins_o[414] = ver_i[284];
  assign ins_o[413] = ver_i[283];
  assign ins_o[412] = ver_i[282];
  assign ins_o[411] = ver_i[281];
  assign ins_o[410] = ver_i[280];
  assign ins_o[409] = ver_i[279];
  assign ins_o[408] = ver_i[278];
  assign ins_o[407] = ver_i[277];
  assign ins_o[406] = ver_i[276];
  assign ins_o[405] = ver_i[275];
  assign ins_o[404] = ver_i[274];
  assign ins_o[403] = ver_i[273];
  assign ins_o[402] = ver_i[272];
  assign ins_o[401] = ver_i[271];
  assign ins_o[400] = ver_i[270];
  assign ins_o[399] = ver_i[269];
  assign ins_o[398] = ver_i[268];
  assign ins_o[397] = ver_i[267];
  assign ins_o[396] = ver_i[266];
  assign ins_o[395] = ver_i[265];
  assign ins_o[394] = ver_i[264];
  assign ins_o[393] = ver_i[263];
  assign ins_o[392] = ver_i[262];
  assign ins_o[391] = ver_i[261];
  assign ins_o[390] = ver_i[260];
  assign ins_o[389] = ver_i[129];
  assign ins_o[388] = ver_i[128];
  assign ins_o[387] = ver_i[127];
  assign ins_o[386] = ver_i[126];
  assign ins_o[385] = ver_i[125];
  assign ins_o[384] = ver_i[124];
  assign ins_o[383] = ver_i[123];
  assign ins_o[382] = ver_i[122];
  assign ins_o[381] = ver_i[121];
  assign ins_o[380] = ver_i[120];
  assign ins_o[379] = ver_i[119];
  assign ins_o[378] = ver_i[118];
  assign ins_o[377] = ver_i[117];
  assign ins_o[376] = ver_i[116];
  assign ins_o[375] = ver_i[115];
  assign ins_o[374] = ver_i[114];
  assign ins_o[373] = ver_i[113];
  assign ins_o[372] = ver_i[112];
  assign ins_o[371] = ver_i[111];
  assign ins_o[370] = ver_i[110];
  assign ins_o[369] = ver_i[109];
  assign ins_o[368] = ver_i[108];
  assign ins_o[367] = ver_i[107];
  assign ins_o[366] = ver_i[106];
  assign ins_o[365] = ver_i[105];
  assign ins_o[364] = ver_i[104];
  assign ins_o[363] = ver_i[103];
  assign ins_o[362] = ver_i[102];
  assign ins_o[361] = ver_i[101];
  assign ins_o[360] = ver_i[100];
  assign ins_o[359] = ver_i[99];
  assign ins_o[358] = ver_i[98];
  assign ins_o[357] = ver_i[97];
  assign ins_o[356] = ver_i[96];
  assign ins_o[355] = ver_i[95];
  assign ins_o[354] = ver_i[94];
  assign ins_o[353] = ver_i[93];
  assign ins_o[352] = ver_i[92];
  assign ins_o[351] = ver_i[91];
  assign ins_o[350] = ver_i[90];
  assign ins_o[349] = ver_i[89];
  assign ins_o[348] = ver_i[88];
  assign ins_o[347] = ver_i[87];
  assign ins_o[346] = ver_i[86];
  assign ins_o[345] = ver_i[85];
  assign ins_o[344] = ver_i[84];
  assign ins_o[343] = ver_i[83];
  assign ins_o[342] = ver_i[82];
  assign ins_o[341] = ver_i[81];
  assign ins_o[340] = ver_i[80];
  assign ins_o[339] = ver_i[79];
  assign ins_o[338] = ver_i[78];
  assign ins_o[337] = ver_i[77];
  assign ins_o[336] = ver_i[76];
  assign ins_o[335] = ver_i[75];
  assign ins_o[334] = ver_i[74];
  assign ins_o[333] = ver_i[73];
  assign ins_o[332] = ver_i[72];
  assign ins_o[331] = ver_i[71];
  assign ins_o[330] = ver_i[70];
  assign ins_o[329] = ver_i[69];
  assign ins_o[328] = ver_i[68];
  assign ins_o[327] = ver_i[67];
  assign ins_o[326] = ver_i[66];
  assign ins_o[325] = ver_i[65];
  assign ins_o[324] = ver_i[64];
  assign ins_o[323] = ver_i[63];
  assign ins_o[322] = ver_i[62];
  assign ins_o[321] = ver_i[61];
  assign ins_o[320] = ver_i[60];
  assign ins_o[319] = ver_i[59];
  assign ins_o[318] = ver_i[58];
  assign ins_o[317] = ver_i[57];
  assign ins_o[316] = ver_i[56];
  assign ins_o[315] = ver_i[55];
  assign ins_o[314] = ver_i[54];
  assign ins_o[313] = ver_i[53];
  assign ins_o[312] = ver_i[52];
  assign ins_o[311] = ver_i[51];
  assign ins_o[310] = ver_i[50];
  assign ins_o[309] = ver_i[49];
  assign ins_o[308] = ver_i[48];
  assign ins_o[307] = ver_i[47];
  assign ins_o[306] = ver_i[46];
  assign ins_o[305] = ver_i[45];
  assign ins_o[304] = ver_i[44];
  assign ins_o[303] = ver_i[43];
  assign ins_o[302] = ver_i[42];
  assign ins_o[301] = ver_i[41];
  assign ins_o[300] = ver_i[40];
  assign ins_o[299] = ver_i[39];
  assign ins_o[298] = ver_i[38];
  assign ins_o[297] = ver_i[37];
  assign ins_o[296] = ver_i[36];
  assign ins_o[295] = ver_i[35];
  assign ins_o[294] = ver_i[34];
  assign ins_o[293] = ver_i[33];
  assign ins_o[292] = ver_i[32];
  assign ins_o[291] = ver_i[31];
  assign ins_o[290] = ver_i[30];
  assign ins_o[289] = ver_i[29];
  assign ins_o[288] = ver_i[28];
  assign ins_o[287] = ver_i[27];
  assign ins_o[286] = ver_i[26];
  assign ins_o[285] = ver_i[25];
  assign ins_o[284] = ver_i[24];
  assign ins_o[283] = ver_i[23];
  assign ins_o[282] = ver_i[22];
  assign ins_o[281] = ver_i[21];
  assign ins_o[280] = ver_i[20];
  assign ins_o[279] = ver_i[19];
  assign ins_o[278] = ver_i[18];
  assign ins_o[277] = ver_i[17];
  assign ins_o[276] = ver_i[16];
  assign ins_o[275] = ver_i[15];
  assign ins_o[274] = ver_i[14];
  assign ins_o[273] = ver_i[13];
  assign ins_o[272] = ver_i[12];
  assign ins_o[271] = ver_i[11];
  assign ins_o[270] = ver_i[10];
  assign ins_o[269] = ver_i[9];
  assign ins_o[268] = ver_i[8];
  assign ins_o[267] = ver_i[7];
  assign ins_o[266] = ver_i[6];
  assign ins_o[265] = ver_i[5];
  assign ins_o[264] = ver_i[4];
  assign ins_o[263] = ver_i[3];
  assign ins_o[262] = ver_i[2];
  assign ins_o[261] = ver_i[1];
  assign ins_o[260] = ver_i[0];
  assign ins_o[259] = outs_i[649];
  assign ins_o[258] = outs_i[648];
  assign ins_o[257] = outs_i[647];
  assign ins_o[256] = outs_i[646];
  assign ins_o[255] = outs_i[645];
  assign ins_o[254] = outs_i[644];
  assign ins_o[253] = outs_i[643];
  assign ins_o[252] = outs_i[642];
  assign ins_o[251] = outs_i[641];
  assign ins_o[250] = outs_i[640];
  assign ins_o[249] = outs_i[639];
  assign ins_o[248] = outs_i[638];
  assign ins_o[247] = outs_i[637];
  assign ins_o[246] = outs_i[636];
  assign ins_o[245] = outs_i[635];
  assign ins_o[244] = outs_i[634];
  assign ins_o[243] = outs_i[633];
  assign ins_o[242] = outs_i[632];
  assign ins_o[241] = outs_i[631];
  assign ins_o[240] = outs_i[630];
  assign ins_o[239] = outs_i[629];
  assign ins_o[238] = outs_i[628];
  assign ins_o[237] = outs_i[627];
  assign ins_o[236] = outs_i[626];
  assign ins_o[235] = outs_i[625];
  assign ins_o[234] = outs_i[624];
  assign ins_o[233] = outs_i[623];
  assign ins_o[232] = outs_i[622];
  assign ins_o[231] = outs_i[621];
  assign ins_o[230] = outs_i[620];
  assign ins_o[229] = outs_i[619];
  assign ins_o[228] = outs_i[618];
  assign ins_o[227] = outs_i[617];
  assign ins_o[226] = outs_i[616];
  assign ins_o[225] = outs_i[615];
  assign ins_o[224] = outs_i[614];
  assign ins_o[223] = outs_i[613];
  assign ins_o[222] = outs_i[612];
  assign ins_o[221] = outs_i[611];
  assign ins_o[220] = outs_i[610];
  assign ins_o[219] = outs_i[609];
  assign ins_o[218] = outs_i[608];
  assign ins_o[217] = outs_i[607];
  assign ins_o[216] = outs_i[606];
  assign ins_o[215] = outs_i[605];
  assign ins_o[214] = outs_i[604];
  assign ins_o[213] = outs_i[603];
  assign ins_o[212] = outs_i[602];
  assign ins_o[211] = outs_i[601];
  assign ins_o[210] = outs_i[600];
  assign ins_o[209] = outs_i[599];
  assign ins_o[208] = outs_i[598];
  assign ins_o[207] = outs_i[597];
  assign ins_o[206] = outs_i[596];
  assign ins_o[205] = outs_i[595];
  assign ins_o[204] = outs_i[594];
  assign ins_o[203] = outs_i[593];
  assign ins_o[202] = outs_i[592];
  assign ins_o[201] = outs_i[591];
  assign ins_o[200] = outs_i[590];
  assign ins_o[199] = outs_i[589];
  assign ins_o[198] = outs_i[588];
  assign ins_o[197] = outs_i[587];
  assign ins_o[196] = outs_i[586];
  assign ins_o[195] = outs_i[585];
  assign ins_o[194] = outs_i[584];
  assign ins_o[193] = outs_i[583];
  assign ins_o[192] = outs_i[582];
  assign ins_o[191] = outs_i[581];
  assign ins_o[190] = outs_i[580];
  assign ins_o[189] = outs_i[579];
  assign ins_o[188] = outs_i[578];
  assign ins_o[187] = outs_i[577];
  assign ins_o[186] = outs_i[576];
  assign ins_o[185] = outs_i[575];
  assign ins_o[184] = outs_i[574];
  assign ins_o[183] = outs_i[573];
  assign ins_o[182] = outs_i[572];
  assign ins_o[181] = outs_i[571];
  assign ins_o[180] = outs_i[570];
  assign ins_o[179] = outs_i[569];
  assign ins_o[178] = outs_i[568];
  assign ins_o[177] = outs_i[567];
  assign ins_o[176] = outs_i[566];
  assign ins_o[175] = outs_i[565];
  assign ins_o[174] = outs_i[564];
  assign ins_o[173] = outs_i[563];
  assign ins_o[172] = outs_i[562];
  assign ins_o[171] = outs_i[561];
  assign ins_o[170] = outs_i[560];
  assign ins_o[169] = outs_i[559];
  assign ins_o[168] = outs_i[558];
  assign ins_o[167] = outs_i[557];
  assign ins_o[166] = outs_i[556];
  assign ins_o[165] = outs_i[555];
  assign ins_o[164] = outs_i[554];
  assign ins_o[163] = outs_i[553];
  assign ins_o[162] = outs_i[552];
  assign ins_o[161] = outs_i[551];
  assign ins_o[160] = outs_i[550];
  assign ins_o[159] = outs_i[549];
  assign ins_o[158] = outs_i[548];
  assign ins_o[157] = outs_i[547];
  assign ins_o[156] = outs_i[546];
  assign ins_o[155] = outs_i[545];
  assign ins_o[154] = outs_i[544];
  assign ins_o[153] = outs_i[543];
  assign ins_o[152] = outs_i[542];
  assign ins_o[151] = outs_i[541];
  assign ins_o[150] = outs_i[540];
  assign ins_o[149] = outs_i[539];
  assign ins_o[148] = outs_i[538];
  assign ins_o[147] = outs_i[537];
  assign ins_o[146] = outs_i[536];
  assign ins_o[145] = outs_i[535];
  assign ins_o[144] = outs_i[534];
  assign ins_o[143] = outs_i[533];
  assign ins_o[142] = outs_i[532];
  assign ins_o[141] = outs_i[531];
  assign ins_o[140] = outs_i[530];
  assign ins_o[139] = outs_i[529];
  assign ins_o[138] = outs_i[528];
  assign ins_o[137] = outs_i[527];
  assign ins_o[136] = outs_i[526];
  assign ins_o[135] = outs_i[525];
  assign ins_o[134] = outs_i[524];
  assign ins_o[133] = outs_i[523];
  assign ins_o[132] = outs_i[522];
  assign ins_o[131] = outs_i[521];
  assign ins_o[130] = outs_i[520];
  assign ins_o[129] = hor_i[129];
  assign ins_o[128] = hor_i[128];
  assign ins_o[127] = hor_i[127];
  assign ins_o[126] = hor_i[126];
  assign ins_o[125] = hor_i[125];
  assign ins_o[124] = hor_i[124];
  assign ins_o[123] = hor_i[123];
  assign ins_o[122] = hor_i[122];
  assign ins_o[121] = hor_i[121];
  assign ins_o[120] = hor_i[120];
  assign ins_o[119] = hor_i[119];
  assign ins_o[118] = hor_i[118];
  assign ins_o[117] = hor_i[117];
  assign ins_o[116] = hor_i[116];
  assign ins_o[115] = hor_i[115];
  assign ins_o[114] = hor_i[114];
  assign ins_o[113] = hor_i[113];
  assign ins_o[112] = hor_i[112];
  assign ins_o[111] = hor_i[111];
  assign ins_o[110] = hor_i[110];
  assign ins_o[109] = hor_i[109];
  assign ins_o[108] = hor_i[108];
  assign ins_o[107] = hor_i[107];
  assign ins_o[106] = hor_i[106];
  assign ins_o[105] = hor_i[105];
  assign ins_o[104] = hor_i[104];
  assign ins_o[103] = hor_i[103];
  assign ins_o[102] = hor_i[102];
  assign ins_o[101] = hor_i[101];
  assign ins_o[100] = hor_i[100];
  assign ins_o[99] = hor_i[99];
  assign ins_o[98] = hor_i[98];
  assign ins_o[97] = hor_i[97];
  assign ins_o[96] = hor_i[96];
  assign ins_o[95] = hor_i[95];
  assign ins_o[94] = hor_i[94];
  assign ins_o[93] = hor_i[93];
  assign ins_o[92] = hor_i[92];
  assign ins_o[91] = hor_i[91];
  assign ins_o[90] = hor_i[90];
  assign ins_o[89] = hor_i[89];
  assign ins_o[88] = hor_i[88];
  assign ins_o[87] = hor_i[87];
  assign ins_o[86] = hor_i[86];
  assign ins_o[85] = hor_i[85];
  assign ins_o[84] = hor_i[84];
  assign ins_o[83] = hor_i[83];
  assign ins_o[82] = hor_i[82];
  assign ins_o[81] = hor_i[81];
  assign ins_o[80] = hor_i[80];
  assign ins_o[79] = hor_i[79];
  assign ins_o[78] = hor_i[78];
  assign ins_o[77] = hor_i[77];
  assign ins_o[76] = hor_i[76];
  assign ins_o[75] = hor_i[75];
  assign ins_o[74] = hor_i[74];
  assign ins_o[73] = hor_i[73];
  assign ins_o[72] = hor_i[72];
  assign ins_o[71] = hor_i[71];
  assign ins_o[70] = hor_i[70];
  assign ins_o[69] = hor_i[69];
  assign ins_o[68] = hor_i[68];
  assign ins_o[67] = hor_i[67];
  assign ins_o[66] = hor_i[66];
  assign ins_o[65] = hor_i[65];
  assign ins_o[64] = hor_i[64];
  assign ins_o[63] = hor_i[63];
  assign ins_o[62] = hor_i[62];
  assign ins_o[61] = hor_i[61];
  assign ins_o[60] = hor_i[60];
  assign ins_o[59] = hor_i[59];
  assign ins_o[58] = hor_i[58];
  assign ins_o[57] = hor_i[57];
  assign ins_o[56] = hor_i[56];
  assign ins_o[55] = hor_i[55];
  assign ins_o[54] = hor_i[54];
  assign ins_o[53] = hor_i[53];
  assign ins_o[52] = hor_i[52];
  assign ins_o[51] = hor_i[51];
  assign ins_o[50] = hor_i[50];
  assign ins_o[49] = hor_i[49];
  assign ins_o[48] = hor_i[48];
  assign ins_o[47] = hor_i[47];
  assign ins_o[46] = hor_i[46];
  assign ins_o[45] = hor_i[45];
  assign ins_o[44] = hor_i[44];
  assign ins_o[43] = hor_i[43];
  assign ins_o[42] = hor_i[42];
  assign ins_o[41] = hor_i[41];
  assign ins_o[40] = hor_i[40];
  assign ins_o[39] = hor_i[39];
  assign ins_o[38] = hor_i[38];
  assign ins_o[37] = hor_i[37];
  assign ins_o[36] = hor_i[36];
  assign ins_o[35] = hor_i[35];
  assign ins_o[34] = hor_i[34];
  assign ins_o[33] = hor_i[33];
  assign ins_o[32] = hor_i[32];
  assign ins_o[31] = hor_i[31];
  assign ins_o[30] = hor_i[30];
  assign ins_o[29] = hor_i[29];
  assign ins_o[28] = hor_i[28];
  assign ins_o[27] = hor_i[27];
  assign ins_o[26] = hor_i[26];
  assign ins_o[25] = hor_i[25];
  assign ins_o[24] = hor_i[24];
  assign ins_o[23] = hor_i[23];
  assign ins_o[22] = hor_i[22];
  assign ins_o[21] = hor_i[21];
  assign ins_o[20] = hor_i[20];
  assign ins_o[19] = hor_i[19];
  assign ins_o[18] = hor_i[18];
  assign ins_o[17] = hor_i[17];
  assign ins_o[16] = hor_i[16];
  assign ins_o[15] = hor_i[15];
  assign ins_o[14] = hor_i[14];
  assign ins_o[13] = hor_i[13];
  assign ins_o[12] = hor_i[12];
  assign ins_o[11] = hor_i[11];
  assign ins_o[10] = hor_i[10];
  assign ins_o[9] = hor_i[9];
  assign ins_o[8] = hor_i[8];
  assign ins_o[7] = hor_i[7];
  assign ins_o[6] = hor_i[6];
  assign ins_o[5] = hor_i[5];
  assign ins_o[4] = hor_i[4];
  assign ins_o[3] = hor_i[3];
  assign ins_o[2] = hor_i[2];
  assign ins_o[1] = hor_i[1];
  assign ins_o[0] = hor_i[0];
  assign hor_o[259] = outs_i[779];
  assign hor_o[258] = outs_i[778];
  assign hor_o[257] = outs_i[777];
  assign hor_o[256] = outs_i[776];
  assign hor_o[255] = outs_i[775];
  assign hor_o[254] = outs_i[774];
  assign hor_o[253] = outs_i[773];
  assign hor_o[252] = outs_i[772];
  assign hor_o[251] = outs_i[771];
  assign hor_o[250] = outs_i[770];
  assign hor_o[249] = outs_i[769];
  assign hor_o[248] = outs_i[768];
  assign hor_o[247] = outs_i[767];
  assign hor_o[246] = outs_i[766];
  assign hor_o[245] = outs_i[765];
  assign hor_o[244] = outs_i[764];
  assign hor_o[243] = outs_i[763];
  assign hor_o[242] = outs_i[762];
  assign hor_o[241] = outs_i[761];
  assign hor_o[240] = outs_i[760];
  assign hor_o[239] = outs_i[759];
  assign hor_o[238] = outs_i[758];
  assign hor_o[237] = outs_i[757];
  assign hor_o[236] = outs_i[756];
  assign hor_o[235] = outs_i[755];
  assign hor_o[234] = outs_i[754];
  assign hor_o[233] = outs_i[753];
  assign hor_o[232] = outs_i[752];
  assign hor_o[231] = outs_i[751];
  assign hor_o[230] = outs_i[750];
  assign hor_o[229] = outs_i[749];
  assign hor_o[228] = outs_i[748];
  assign hor_o[227] = outs_i[747];
  assign hor_o[226] = outs_i[746];
  assign hor_o[225] = outs_i[745];
  assign hor_o[224] = outs_i[744];
  assign hor_o[223] = outs_i[743];
  assign hor_o[222] = outs_i[742];
  assign hor_o[221] = outs_i[741];
  assign hor_o[220] = outs_i[740];
  assign hor_o[219] = outs_i[739];
  assign hor_o[218] = outs_i[738];
  assign hor_o[217] = outs_i[737];
  assign hor_o[216] = outs_i[736];
  assign hor_o[215] = outs_i[735];
  assign hor_o[214] = outs_i[734];
  assign hor_o[213] = outs_i[733];
  assign hor_o[212] = outs_i[732];
  assign hor_o[211] = outs_i[731];
  assign hor_o[210] = outs_i[730];
  assign hor_o[209] = outs_i[729];
  assign hor_o[208] = outs_i[728];
  assign hor_o[207] = outs_i[727];
  assign hor_o[206] = outs_i[726];
  assign hor_o[205] = outs_i[725];
  assign hor_o[204] = outs_i[724];
  assign hor_o[203] = outs_i[723];
  assign hor_o[202] = outs_i[722];
  assign hor_o[201] = outs_i[721];
  assign hor_o[200] = outs_i[720];
  assign hor_o[199] = outs_i[719];
  assign hor_o[198] = outs_i[718];
  assign hor_o[197] = outs_i[717];
  assign hor_o[196] = outs_i[716];
  assign hor_o[195] = outs_i[715];
  assign hor_o[194] = outs_i[714];
  assign hor_o[193] = outs_i[713];
  assign hor_o[192] = outs_i[712];
  assign hor_o[191] = outs_i[711];
  assign hor_o[190] = outs_i[710];
  assign hor_o[189] = outs_i[709];
  assign hor_o[188] = outs_i[708];
  assign hor_o[187] = outs_i[707];
  assign hor_o[186] = outs_i[706];
  assign hor_o[185] = outs_i[705];
  assign hor_o[184] = outs_i[704];
  assign hor_o[183] = outs_i[703];
  assign hor_o[182] = outs_i[702];
  assign hor_o[181] = outs_i[701];
  assign hor_o[180] = outs_i[700];
  assign hor_o[179] = outs_i[699];
  assign hor_o[178] = outs_i[698];
  assign hor_o[177] = outs_i[697];
  assign hor_o[176] = outs_i[696];
  assign hor_o[175] = outs_i[695];
  assign hor_o[174] = outs_i[694];
  assign hor_o[173] = outs_i[693];
  assign hor_o[172] = outs_i[692];
  assign hor_o[171] = outs_i[691];
  assign hor_o[170] = outs_i[690];
  assign hor_o[169] = outs_i[689];
  assign hor_o[168] = outs_i[688];
  assign hor_o[167] = outs_i[687];
  assign hor_o[166] = outs_i[686];
  assign hor_o[165] = outs_i[685];
  assign hor_o[164] = outs_i[684];
  assign hor_o[163] = outs_i[683];
  assign hor_o[162] = outs_i[682];
  assign hor_o[161] = outs_i[681];
  assign hor_o[160] = outs_i[680];
  assign hor_o[159] = outs_i[679];
  assign hor_o[158] = outs_i[678];
  assign hor_o[157] = outs_i[677];
  assign hor_o[156] = outs_i[676];
  assign hor_o[155] = outs_i[675];
  assign hor_o[154] = outs_i[674];
  assign hor_o[153] = outs_i[673];
  assign hor_o[152] = outs_i[672];
  assign hor_o[151] = outs_i[671];
  assign hor_o[150] = outs_i[670];
  assign hor_o[149] = outs_i[669];
  assign hor_o[148] = outs_i[668];
  assign hor_o[147] = outs_i[667];
  assign hor_o[146] = outs_i[666];
  assign hor_o[145] = outs_i[665];
  assign hor_o[144] = outs_i[664];
  assign hor_o[143] = outs_i[663];
  assign hor_o[142] = outs_i[662];
  assign hor_o[141] = outs_i[661];
  assign hor_o[140] = outs_i[660];
  assign hor_o[139] = outs_i[659];
  assign hor_o[138] = outs_i[658];
  assign hor_o[137] = outs_i[657];
  assign hor_o[136] = outs_i[656];
  assign hor_o[135] = outs_i[655];
  assign hor_o[134] = outs_i[654];
  assign hor_o[133] = outs_i[653];
  assign hor_o[132] = outs_i[652];
  assign hor_o[131] = outs_i[651];
  assign hor_o[130] = outs_i[650];
  assign hor_o[129] = outs_i[129];
  assign hor_o[128] = outs_i[128];
  assign hor_o[127] = outs_i[127];
  assign hor_o[126] = outs_i[126];
  assign hor_o[125] = outs_i[125];
  assign hor_o[124] = outs_i[124];
  assign hor_o[123] = outs_i[123];
  assign hor_o[122] = outs_i[122];
  assign hor_o[121] = outs_i[121];
  assign hor_o[120] = outs_i[120];
  assign hor_o[119] = outs_i[119];
  assign hor_o[118] = outs_i[118];
  assign hor_o[117] = outs_i[117];
  assign hor_o[116] = outs_i[116];
  assign hor_o[115] = outs_i[115];
  assign hor_o[114] = outs_i[114];
  assign hor_o[113] = outs_i[113];
  assign hor_o[112] = outs_i[112];
  assign hor_o[111] = outs_i[111];
  assign hor_o[110] = outs_i[110];
  assign hor_o[109] = outs_i[109];
  assign hor_o[108] = outs_i[108];
  assign hor_o[107] = outs_i[107];
  assign hor_o[106] = outs_i[106];
  assign hor_o[105] = outs_i[105];
  assign hor_o[104] = outs_i[104];
  assign hor_o[103] = outs_i[103];
  assign hor_o[102] = outs_i[102];
  assign hor_o[101] = outs_i[101];
  assign hor_o[100] = outs_i[100];
  assign hor_o[99] = outs_i[99];
  assign hor_o[98] = outs_i[98];
  assign hor_o[97] = outs_i[97];
  assign hor_o[96] = outs_i[96];
  assign hor_o[95] = outs_i[95];
  assign hor_o[94] = outs_i[94];
  assign hor_o[93] = outs_i[93];
  assign hor_o[92] = outs_i[92];
  assign hor_o[91] = outs_i[91];
  assign hor_o[90] = outs_i[90];
  assign hor_o[89] = outs_i[89];
  assign hor_o[88] = outs_i[88];
  assign hor_o[87] = outs_i[87];
  assign hor_o[86] = outs_i[86];
  assign hor_o[85] = outs_i[85];
  assign hor_o[84] = outs_i[84];
  assign hor_o[83] = outs_i[83];
  assign hor_o[82] = outs_i[82];
  assign hor_o[81] = outs_i[81];
  assign hor_o[80] = outs_i[80];
  assign hor_o[79] = outs_i[79];
  assign hor_o[78] = outs_i[78];
  assign hor_o[77] = outs_i[77];
  assign hor_o[76] = outs_i[76];
  assign hor_o[75] = outs_i[75];
  assign hor_o[74] = outs_i[74];
  assign hor_o[73] = outs_i[73];
  assign hor_o[72] = outs_i[72];
  assign hor_o[71] = outs_i[71];
  assign hor_o[70] = outs_i[70];
  assign hor_o[69] = outs_i[69];
  assign hor_o[68] = outs_i[68];
  assign hor_o[67] = outs_i[67];
  assign hor_o[66] = outs_i[66];
  assign hor_o[65] = outs_i[65];
  assign hor_o[64] = outs_i[64];
  assign hor_o[63] = outs_i[63];
  assign hor_o[62] = outs_i[62];
  assign hor_o[61] = outs_i[61];
  assign hor_o[60] = outs_i[60];
  assign hor_o[59] = outs_i[59];
  assign hor_o[58] = outs_i[58];
  assign hor_o[57] = outs_i[57];
  assign hor_o[56] = outs_i[56];
  assign hor_o[55] = outs_i[55];
  assign hor_o[54] = outs_i[54];
  assign hor_o[53] = outs_i[53];
  assign hor_o[52] = outs_i[52];
  assign hor_o[51] = outs_i[51];
  assign hor_o[50] = outs_i[50];
  assign hor_o[49] = outs_i[49];
  assign hor_o[48] = outs_i[48];
  assign hor_o[47] = outs_i[47];
  assign hor_o[46] = outs_i[46];
  assign hor_o[45] = outs_i[45];
  assign hor_o[44] = outs_i[44];
  assign hor_o[43] = outs_i[43];
  assign hor_o[42] = outs_i[42];
  assign hor_o[41] = outs_i[41];
  assign hor_o[40] = outs_i[40];
  assign hor_o[39] = outs_i[39];
  assign hor_o[38] = outs_i[38];
  assign hor_o[37] = outs_i[37];
  assign hor_o[36] = outs_i[36];
  assign hor_o[35] = outs_i[35];
  assign hor_o[34] = outs_i[34];
  assign hor_o[33] = outs_i[33];
  assign hor_o[32] = outs_i[32];
  assign hor_o[31] = outs_i[31];
  assign hor_o[30] = outs_i[30];
  assign hor_o[29] = outs_i[29];
  assign hor_o[28] = outs_i[28];
  assign hor_o[27] = outs_i[27];
  assign hor_o[26] = outs_i[26];
  assign hor_o[25] = outs_i[25];
  assign hor_o[24] = outs_i[24];
  assign hor_o[23] = outs_i[23];
  assign hor_o[22] = outs_i[22];
  assign hor_o[21] = outs_i[21];
  assign hor_o[20] = outs_i[20];
  assign hor_o[19] = outs_i[19];
  assign hor_o[18] = outs_i[18];
  assign hor_o[17] = outs_i[17];
  assign hor_o[16] = outs_i[16];
  assign hor_o[15] = outs_i[15];
  assign hor_o[14] = outs_i[14];
  assign hor_o[13] = outs_i[13];
  assign hor_o[12] = outs_i[12];
  assign hor_o[11] = outs_i[11];
  assign hor_o[10] = outs_i[10];
  assign hor_o[9] = outs_i[9];
  assign hor_o[8] = outs_i[8];
  assign hor_o[7] = outs_i[7];
  assign hor_o[6] = outs_i[6];
  assign hor_o[5] = outs_i[5];
  assign hor_o[4] = outs_i[4];
  assign hor_o[3] = outs_i[3];
  assign hor_o[2] = outs_i[2];
  assign hor_o[1] = outs_i[1];
  assign hor_o[0] = outs_i[0];
  assign ver_o[519] = outs_i[1039];
  assign ver_o[518] = outs_i[1038];
  assign ver_o[517] = outs_i[1037];
  assign ver_o[516] = outs_i[1036];
  assign ver_o[515] = outs_i[1035];
  assign ver_o[514] = outs_i[1034];
  assign ver_o[513] = outs_i[1033];
  assign ver_o[512] = outs_i[1032];
  assign ver_o[511] = outs_i[1031];
  assign ver_o[510] = outs_i[1030];
  assign ver_o[509] = outs_i[1029];
  assign ver_o[508] = outs_i[1028];
  assign ver_o[507] = outs_i[1027];
  assign ver_o[506] = outs_i[1026];
  assign ver_o[505] = outs_i[1025];
  assign ver_o[504] = outs_i[1024];
  assign ver_o[503] = outs_i[1023];
  assign ver_o[502] = outs_i[1022];
  assign ver_o[501] = outs_i[1021];
  assign ver_o[500] = outs_i[1020];
  assign ver_o[499] = outs_i[1019];
  assign ver_o[498] = outs_i[1018];
  assign ver_o[497] = outs_i[1017];
  assign ver_o[496] = outs_i[1016];
  assign ver_o[495] = outs_i[1015];
  assign ver_o[494] = outs_i[1014];
  assign ver_o[493] = outs_i[1013];
  assign ver_o[492] = outs_i[1012];
  assign ver_o[491] = outs_i[1011];
  assign ver_o[490] = outs_i[1010];
  assign ver_o[489] = outs_i[1009];
  assign ver_o[488] = outs_i[1008];
  assign ver_o[487] = outs_i[1007];
  assign ver_o[486] = outs_i[1006];
  assign ver_o[485] = outs_i[1005];
  assign ver_o[484] = outs_i[1004];
  assign ver_o[483] = outs_i[1003];
  assign ver_o[482] = outs_i[1002];
  assign ver_o[481] = outs_i[1001];
  assign ver_o[480] = outs_i[1000];
  assign ver_o[479] = outs_i[999];
  assign ver_o[478] = outs_i[998];
  assign ver_o[477] = outs_i[997];
  assign ver_o[476] = outs_i[996];
  assign ver_o[475] = outs_i[995];
  assign ver_o[474] = outs_i[994];
  assign ver_o[473] = outs_i[993];
  assign ver_o[472] = outs_i[992];
  assign ver_o[471] = outs_i[991];
  assign ver_o[470] = outs_i[990];
  assign ver_o[469] = outs_i[989];
  assign ver_o[468] = outs_i[988];
  assign ver_o[467] = outs_i[987];
  assign ver_o[466] = outs_i[986];
  assign ver_o[465] = outs_i[985];
  assign ver_o[464] = outs_i[984];
  assign ver_o[463] = outs_i[983];
  assign ver_o[462] = outs_i[982];
  assign ver_o[461] = outs_i[981];
  assign ver_o[460] = outs_i[980];
  assign ver_o[459] = outs_i[979];
  assign ver_o[458] = outs_i[978];
  assign ver_o[457] = outs_i[977];
  assign ver_o[456] = outs_i[976];
  assign ver_o[455] = outs_i[975];
  assign ver_o[454] = outs_i[974];
  assign ver_o[453] = outs_i[973];
  assign ver_o[452] = outs_i[972];
  assign ver_o[451] = outs_i[971];
  assign ver_o[450] = outs_i[970];
  assign ver_o[449] = outs_i[969];
  assign ver_o[448] = outs_i[968];
  assign ver_o[447] = outs_i[967];
  assign ver_o[446] = outs_i[966];
  assign ver_o[445] = outs_i[965];
  assign ver_o[444] = outs_i[964];
  assign ver_o[443] = outs_i[963];
  assign ver_o[442] = outs_i[962];
  assign ver_o[441] = outs_i[961];
  assign ver_o[440] = outs_i[960];
  assign ver_o[439] = outs_i[959];
  assign ver_o[438] = outs_i[958];
  assign ver_o[437] = outs_i[957];
  assign ver_o[436] = outs_i[956];
  assign ver_o[435] = outs_i[955];
  assign ver_o[434] = outs_i[954];
  assign ver_o[433] = outs_i[953];
  assign ver_o[432] = outs_i[952];
  assign ver_o[431] = outs_i[951];
  assign ver_o[430] = outs_i[950];
  assign ver_o[429] = outs_i[949];
  assign ver_o[428] = outs_i[948];
  assign ver_o[427] = outs_i[947];
  assign ver_o[426] = outs_i[946];
  assign ver_o[425] = outs_i[945];
  assign ver_o[424] = outs_i[944];
  assign ver_o[423] = outs_i[943];
  assign ver_o[422] = outs_i[942];
  assign ver_o[421] = outs_i[941];
  assign ver_o[420] = outs_i[940];
  assign ver_o[419] = outs_i[939];
  assign ver_o[418] = outs_i[938];
  assign ver_o[417] = outs_i[937];
  assign ver_o[416] = outs_i[936];
  assign ver_o[415] = outs_i[935];
  assign ver_o[414] = outs_i[934];
  assign ver_o[413] = outs_i[933];
  assign ver_o[412] = outs_i[932];
  assign ver_o[411] = outs_i[931];
  assign ver_o[410] = outs_i[930];
  assign ver_o[409] = outs_i[929];
  assign ver_o[408] = outs_i[928];
  assign ver_o[407] = outs_i[927];
  assign ver_o[406] = outs_i[926];
  assign ver_o[405] = outs_i[925];
  assign ver_o[404] = outs_i[924];
  assign ver_o[403] = outs_i[923];
  assign ver_o[402] = outs_i[922];
  assign ver_o[401] = outs_i[921];
  assign ver_o[400] = outs_i[920];
  assign ver_o[399] = outs_i[919];
  assign ver_o[398] = outs_i[918];
  assign ver_o[397] = outs_i[917];
  assign ver_o[396] = outs_i[916];
  assign ver_o[395] = outs_i[915];
  assign ver_o[394] = outs_i[914];
  assign ver_o[393] = outs_i[913];
  assign ver_o[392] = outs_i[912];
  assign ver_o[391] = outs_i[911];
  assign ver_o[390] = outs_i[910];
  assign ver_o[389] = outs_i[519];
  assign ver_o[388] = outs_i[518];
  assign ver_o[387] = outs_i[517];
  assign ver_o[386] = outs_i[516];
  assign ver_o[385] = outs_i[515];
  assign ver_o[384] = outs_i[514];
  assign ver_o[383] = outs_i[513];
  assign ver_o[382] = outs_i[512];
  assign ver_o[381] = outs_i[511];
  assign ver_o[380] = outs_i[510];
  assign ver_o[379] = outs_i[509];
  assign ver_o[378] = outs_i[508];
  assign ver_o[377] = outs_i[507];
  assign ver_o[376] = outs_i[506];
  assign ver_o[375] = outs_i[505];
  assign ver_o[374] = outs_i[504];
  assign ver_o[373] = outs_i[503];
  assign ver_o[372] = outs_i[502];
  assign ver_o[371] = outs_i[501];
  assign ver_o[370] = outs_i[500];
  assign ver_o[369] = outs_i[499];
  assign ver_o[368] = outs_i[498];
  assign ver_o[367] = outs_i[497];
  assign ver_o[366] = outs_i[496];
  assign ver_o[365] = outs_i[495];
  assign ver_o[364] = outs_i[494];
  assign ver_o[363] = outs_i[493];
  assign ver_o[362] = outs_i[492];
  assign ver_o[361] = outs_i[491];
  assign ver_o[360] = outs_i[490];
  assign ver_o[359] = outs_i[489];
  assign ver_o[358] = outs_i[488];
  assign ver_o[357] = outs_i[487];
  assign ver_o[356] = outs_i[486];
  assign ver_o[355] = outs_i[485];
  assign ver_o[354] = outs_i[484];
  assign ver_o[353] = outs_i[483];
  assign ver_o[352] = outs_i[482];
  assign ver_o[351] = outs_i[481];
  assign ver_o[350] = outs_i[480];
  assign ver_o[349] = outs_i[479];
  assign ver_o[348] = outs_i[478];
  assign ver_o[347] = outs_i[477];
  assign ver_o[346] = outs_i[476];
  assign ver_o[345] = outs_i[475];
  assign ver_o[344] = outs_i[474];
  assign ver_o[343] = outs_i[473];
  assign ver_o[342] = outs_i[472];
  assign ver_o[341] = outs_i[471];
  assign ver_o[340] = outs_i[470];
  assign ver_o[339] = outs_i[469];
  assign ver_o[338] = outs_i[468];
  assign ver_o[337] = outs_i[467];
  assign ver_o[336] = outs_i[466];
  assign ver_o[335] = outs_i[465];
  assign ver_o[334] = outs_i[464];
  assign ver_o[333] = outs_i[463];
  assign ver_o[332] = outs_i[462];
  assign ver_o[331] = outs_i[461];
  assign ver_o[330] = outs_i[460];
  assign ver_o[329] = outs_i[459];
  assign ver_o[328] = outs_i[458];
  assign ver_o[327] = outs_i[457];
  assign ver_o[326] = outs_i[456];
  assign ver_o[325] = outs_i[455];
  assign ver_o[324] = outs_i[454];
  assign ver_o[323] = outs_i[453];
  assign ver_o[322] = outs_i[452];
  assign ver_o[321] = outs_i[451];
  assign ver_o[320] = outs_i[450];
  assign ver_o[319] = outs_i[449];
  assign ver_o[318] = outs_i[448];
  assign ver_o[317] = outs_i[447];
  assign ver_o[316] = outs_i[446];
  assign ver_o[315] = outs_i[445];
  assign ver_o[314] = outs_i[444];
  assign ver_o[313] = outs_i[443];
  assign ver_o[312] = outs_i[442];
  assign ver_o[311] = outs_i[441];
  assign ver_o[310] = outs_i[440];
  assign ver_o[309] = outs_i[439];
  assign ver_o[308] = outs_i[438];
  assign ver_o[307] = outs_i[437];
  assign ver_o[306] = outs_i[436];
  assign ver_o[305] = outs_i[435];
  assign ver_o[304] = outs_i[434];
  assign ver_o[303] = outs_i[433];
  assign ver_o[302] = outs_i[432];
  assign ver_o[301] = outs_i[431];
  assign ver_o[300] = outs_i[430];
  assign ver_o[299] = outs_i[429];
  assign ver_o[298] = outs_i[428];
  assign ver_o[297] = outs_i[427];
  assign ver_o[296] = outs_i[426];
  assign ver_o[295] = outs_i[425];
  assign ver_o[294] = outs_i[424];
  assign ver_o[293] = outs_i[423];
  assign ver_o[292] = outs_i[422];
  assign ver_o[291] = outs_i[421];
  assign ver_o[290] = outs_i[420];
  assign ver_o[289] = outs_i[419];
  assign ver_o[288] = outs_i[418];
  assign ver_o[287] = outs_i[417];
  assign ver_o[286] = outs_i[416];
  assign ver_o[285] = outs_i[415];
  assign ver_o[284] = outs_i[414];
  assign ver_o[283] = outs_i[413];
  assign ver_o[282] = outs_i[412];
  assign ver_o[281] = outs_i[411];
  assign ver_o[280] = outs_i[410];
  assign ver_o[279] = outs_i[409];
  assign ver_o[278] = outs_i[408];
  assign ver_o[277] = outs_i[407];
  assign ver_o[276] = outs_i[406];
  assign ver_o[275] = outs_i[405];
  assign ver_o[274] = outs_i[404];
  assign ver_o[273] = outs_i[403];
  assign ver_o[272] = outs_i[402];
  assign ver_o[271] = outs_i[401];
  assign ver_o[270] = outs_i[400];
  assign ver_o[269] = outs_i[399];
  assign ver_o[268] = outs_i[398];
  assign ver_o[267] = outs_i[397];
  assign ver_o[266] = outs_i[396];
  assign ver_o[265] = outs_i[395];
  assign ver_o[264] = outs_i[394];
  assign ver_o[263] = outs_i[393];
  assign ver_o[262] = outs_i[392];
  assign ver_o[261] = outs_i[391];
  assign ver_o[260] = outs_i[390];
  assign ver_o[259] = outs_i[909];
  assign ver_o[258] = outs_i[908];
  assign ver_o[257] = outs_i[907];
  assign ver_o[256] = outs_i[906];
  assign ver_o[255] = outs_i[905];
  assign ver_o[254] = outs_i[904];
  assign ver_o[253] = outs_i[903];
  assign ver_o[252] = outs_i[902];
  assign ver_o[251] = outs_i[901];
  assign ver_o[250] = outs_i[900];
  assign ver_o[249] = outs_i[899];
  assign ver_o[248] = outs_i[898];
  assign ver_o[247] = outs_i[897];
  assign ver_o[246] = outs_i[896];
  assign ver_o[245] = outs_i[895];
  assign ver_o[244] = outs_i[894];
  assign ver_o[243] = outs_i[893];
  assign ver_o[242] = outs_i[892];
  assign ver_o[241] = outs_i[891];
  assign ver_o[240] = outs_i[890];
  assign ver_o[239] = outs_i[889];
  assign ver_o[238] = outs_i[888];
  assign ver_o[237] = outs_i[887];
  assign ver_o[236] = outs_i[886];
  assign ver_o[235] = outs_i[885];
  assign ver_o[234] = outs_i[884];
  assign ver_o[233] = outs_i[883];
  assign ver_o[232] = outs_i[882];
  assign ver_o[231] = outs_i[881];
  assign ver_o[230] = outs_i[880];
  assign ver_o[229] = outs_i[879];
  assign ver_o[228] = outs_i[878];
  assign ver_o[227] = outs_i[877];
  assign ver_o[226] = outs_i[876];
  assign ver_o[225] = outs_i[875];
  assign ver_o[224] = outs_i[874];
  assign ver_o[223] = outs_i[873];
  assign ver_o[222] = outs_i[872];
  assign ver_o[221] = outs_i[871];
  assign ver_o[220] = outs_i[870];
  assign ver_o[219] = outs_i[869];
  assign ver_o[218] = outs_i[868];
  assign ver_o[217] = outs_i[867];
  assign ver_o[216] = outs_i[866];
  assign ver_o[215] = outs_i[865];
  assign ver_o[214] = outs_i[864];
  assign ver_o[213] = outs_i[863];
  assign ver_o[212] = outs_i[862];
  assign ver_o[211] = outs_i[861];
  assign ver_o[210] = outs_i[860];
  assign ver_o[209] = outs_i[859];
  assign ver_o[208] = outs_i[858];
  assign ver_o[207] = outs_i[857];
  assign ver_o[206] = outs_i[856];
  assign ver_o[205] = outs_i[855];
  assign ver_o[204] = outs_i[854];
  assign ver_o[203] = outs_i[853];
  assign ver_o[202] = outs_i[852];
  assign ver_o[201] = outs_i[851];
  assign ver_o[200] = outs_i[850];
  assign ver_o[199] = outs_i[849];
  assign ver_o[198] = outs_i[848];
  assign ver_o[197] = outs_i[847];
  assign ver_o[196] = outs_i[846];
  assign ver_o[195] = outs_i[845];
  assign ver_o[194] = outs_i[844];
  assign ver_o[193] = outs_i[843];
  assign ver_o[192] = outs_i[842];
  assign ver_o[191] = outs_i[841];
  assign ver_o[190] = outs_i[840];
  assign ver_o[189] = outs_i[839];
  assign ver_o[188] = outs_i[838];
  assign ver_o[187] = outs_i[837];
  assign ver_o[186] = outs_i[836];
  assign ver_o[185] = outs_i[835];
  assign ver_o[184] = outs_i[834];
  assign ver_o[183] = outs_i[833];
  assign ver_o[182] = outs_i[832];
  assign ver_o[181] = outs_i[831];
  assign ver_o[180] = outs_i[830];
  assign ver_o[179] = outs_i[829];
  assign ver_o[178] = outs_i[828];
  assign ver_o[177] = outs_i[827];
  assign ver_o[176] = outs_i[826];
  assign ver_o[175] = outs_i[825];
  assign ver_o[174] = outs_i[824];
  assign ver_o[173] = outs_i[823];
  assign ver_o[172] = outs_i[822];
  assign ver_o[171] = outs_i[821];
  assign ver_o[170] = outs_i[820];
  assign ver_o[169] = outs_i[819];
  assign ver_o[168] = outs_i[818];
  assign ver_o[167] = outs_i[817];
  assign ver_o[166] = outs_i[816];
  assign ver_o[165] = outs_i[815];
  assign ver_o[164] = outs_i[814];
  assign ver_o[163] = outs_i[813];
  assign ver_o[162] = outs_i[812];
  assign ver_o[161] = outs_i[811];
  assign ver_o[160] = outs_i[810];
  assign ver_o[159] = outs_i[809];
  assign ver_o[158] = outs_i[808];
  assign ver_o[157] = outs_i[807];
  assign ver_o[156] = outs_i[806];
  assign ver_o[155] = outs_i[805];
  assign ver_o[154] = outs_i[804];
  assign ver_o[153] = outs_i[803];
  assign ver_o[152] = outs_i[802];
  assign ver_o[151] = outs_i[801];
  assign ver_o[150] = outs_i[800];
  assign ver_o[149] = outs_i[799];
  assign ver_o[148] = outs_i[798];
  assign ver_o[147] = outs_i[797];
  assign ver_o[146] = outs_i[796];
  assign ver_o[145] = outs_i[795];
  assign ver_o[144] = outs_i[794];
  assign ver_o[143] = outs_i[793];
  assign ver_o[142] = outs_i[792];
  assign ver_o[141] = outs_i[791];
  assign ver_o[140] = outs_i[790];
  assign ver_o[139] = outs_i[789];
  assign ver_o[138] = outs_i[788];
  assign ver_o[137] = outs_i[787];
  assign ver_o[136] = outs_i[786];
  assign ver_o[135] = outs_i[785];
  assign ver_o[134] = outs_i[784];
  assign ver_o[133] = outs_i[783];
  assign ver_o[132] = outs_i[782];
  assign ver_o[131] = outs_i[781];
  assign ver_o[130] = outs_i[780];
  assign ver_o[129] = outs_i[389];
  assign ver_o[128] = outs_i[388];
  assign ver_o[127] = outs_i[387];
  assign ver_o[126] = outs_i[386];
  assign ver_o[125] = outs_i[385];
  assign ver_o[124] = outs_i[384];
  assign ver_o[123] = outs_i[383];
  assign ver_o[122] = outs_i[382];
  assign ver_o[121] = outs_i[381];
  assign ver_o[120] = outs_i[380];
  assign ver_o[119] = outs_i[379];
  assign ver_o[118] = outs_i[378];
  assign ver_o[117] = outs_i[377];
  assign ver_o[116] = outs_i[376];
  assign ver_o[115] = outs_i[375];
  assign ver_o[114] = outs_i[374];
  assign ver_o[113] = outs_i[373];
  assign ver_o[112] = outs_i[372];
  assign ver_o[111] = outs_i[371];
  assign ver_o[110] = outs_i[370];
  assign ver_o[109] = outs_i[369];
  assign ver_o[108] = outs_i[368];
  assign ver_o[107] = outs_i[367];
  assign ver_o[106] = outs_i[366];
  assign ver_o[105] = outs_i[365];
  assign ver_o[104] = outs_i[364];
  assign ver_o[103] = outs_i[363];
  assign ver_o[102] = outs_i[362];
  assign ver_o[101] = outs_i[361];
  assign ver_o[100] = outs_i[360];
  assign ver_o[99] = outs_i[359];
  assign ver_o[98] = outs_i[358];
  assign ver_o[97] = outs_i[357];
  assign ver_o[96] = outs_i[356];
  assign ver_o[95] = outs_i[355];
  assign ver_o[94] = outs_i[354];
  assign ver_o[93] = outs_i[353];
  assign ver_o[92] = outs_i[352];
  assign ver_o[91] = outs_i[351];
  assign ver_o[90] = outs_i[350];
  assign ver_o[89] = outs_i[349];
  assign ver_o[88] = outs_i[348];
  assign ver_o[87] = outs_i[347];
  assign ver_o[86] = outs_i[346];
  assign ver_o[85] = outs_i[345];
  assign ver_o[84] = outs_i[344];
  assign ver_o[83] = outs_i[343];
  assign ver_o[82] = outs_i[342];
  assign ver_o[81] = outs_i[341];
  assign ver_o[80] = outs_i[340];
  assign ver_o[79] = outs_i[339];
  assign ver_o[78] = outs_i[338];
  assign ver_o[77] = outs_i[337];
  assign ver_o[76] = outs_i[336];
  assign ver_o[75] = outs_i[335];
  assign ver_o[74] = outs_i[334];
  assign ver_o[73] = outs_i[333];
  assign ver_o[72] = outs_i[332];
  assign ver_o[71] = outs_i[331];
  assign ver_o[70] = outs_i[330];
  assign ver_o[69] = outs_i[329];
  assign ver_o[68] = outs_i[328];
  assign ver_o[67] = outs_i[327];
  assign ver_o[66] = outs_i[326];
  assign ver_o[65] = outs_i[325];
  assign ver_o[64] = outs_i[324];
  assign ver_o[63] = outs_i[323];
  assign ver_o[62] = outs_i[322];
  assign ver_o[61] = outs_i[321];
  assign ver_o[60] = outs_i[320];
  assign ver_o[59] = outs_i[319];
  assign ver_o[58] = outs_i[318];
  assign ver_o[57] = outs_i[317];
  assign ver_o[56] = outs_i[316];
  assign ver_o[55] = outs_i[315];
  assign ver_o[54] = outs_i[314];
  assign ver_o[53] = outs_i[313];
  assign ver_o[52] = outs_i[312];
  assign ver_o[51] = outs_i[311];
  assign ver_o[50] = outs_i[310];
  assign ver_o[49] = outs_i[309];
  assign ver_o[48] = outs_i[308];
  assign ver_o[47] = outs_i[307];
  assign ver_o[46] = outs_i[306];
  assign ver_o[45] = outs_i[305];
  assign ver_o[44] = outs_i[304];
  assign ver_o[43] = outs_i[303];
  assign ver_o[42] = outs_i[302];
  assign ver_o[41] = outs_i[301];
  assign ver_o[40] = outs_i[300];
  assign ver_o[39] = outs_i[299];
  assign ver_o[38] = outs_i[298];
  assign ver_o[37] = outs_i[297];
  assign ver_o[36] = outs_i[296];
  assign ver_o[35] = outs_i[295];
  assign ver_o[34] = outs_i[294];
  assign ver_o[33] = outs_i[293];
  assign ver_o[32] = outs_i[292];
  assign ver_o[31] = outs_i[291];
  assign ver_o[30] = outs_i[290];
  assign ver_o[29] = outs_i[289];
  assign ver_o[28] = outs_i[288];
  assign ver_o[27] = outs_i[287];
  assign ver_o[26] = outs_i[286];
  assign ver_o[25] = outs_i[285];
  assign ver_o[24] = outs_i[284];
  assign ver_o[23] = outs_i[283];
  assign ver_o[22] = outs_i[282];
  assign ver_o[21] = outs_i[281];
  assign ver_o[20] = outs_i[280];
  assign ver_o[19] = outs_i[279];
  assign ver_o[18] = outs_i[278];
  assign ver_o[17] = outs_i[277];
  assign ver_o[16] = outs_i[276];
  assign ver_o[15] = outs_i[275];
  assign ver_o[14] = outs_i[274];
  assign ver_o[13] = outs_i[273];
  assign ver_o[12] = outs_i[272];
  assign ver_o[11] = outs_i[271];
  assign ver_o[10] = outs_i[270];
  assign ver_o[9] = outs_i[269];
  assign ver_o[8] = outs_i[268];
  assign ver_o[7] = outs_i[267];
  assign ver_o[6] = outs_i[266];
  assign ver_o[5] = outs_i[265];
  assign ver_o[4] = outs_i[264];
  assign ver_o[3] = outs_i[263];
  assign ver_o[2] = outs_i[262];
  assign ver_o[1] = outs_i[261];
  assign ver_o[0] = outs_i[260];

endmodule

